library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity register3 is
    Port ( clk : in  STD_LOGIC;
			  rst : in STD_LOGIC;
           input : in  STD_LOGIC_VECTOR (2 downto 0);
           writeEnable : in  STD_LOGIC;
           output : out  STD_LOGIC_VECTOR (2 downto 0));
end register3;

architecture Behavioral of register3 is
signal tempOut : STD_LOGIC_VECTOR (2 downto 0);

begin
	process (clk, rst) 
	begin
		if (rising_edge(clk)) then
			if (rst = '1') then 
				tempOut <= (others => '0');
			elsif (writeEnable = '1') then 
				tempOut <= input;
			end if;
		end if;
	end process;
	
	output <= tempOut after 10ns;
end Behavioral;

--add testbentch for both registers

